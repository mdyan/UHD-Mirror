//
// Copyright 2011 Ettus Research LLC
//
// This program is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <http://www.gnu.org/licenses/>.
//


// Triple fifo mux (0,1,2)... fair sharing only.

module fifo36_three_way
  #(parameter prio = 1'b0)
   (input clk, input reset, input clear,
    input [35:0] data0_i, input src0_rdy_i, output dst0_rdy_o,
    input [35:0] data1_i, input src1_rdy_i, output dst1_rdy_o,
    input [35:0] data2_i, input src2_rdy_i, output dst2_rdy_o,
    output [35:0] data_o, output src_rdy_o, input dst_rdy_i);

   wire [35:0] 	  data0_int, data1_int, data2_int;
   wire 	  src0_rdy_int, dst0_rdy_int, src1_rdy_int, dst1_rdy_int, src2_rdy_int, dst2_rdy_int;
   
   fifo_short #(.WIDTH(36)) mux_fifo_in0
     (.clk(clk), .reset(reset), .clear(clear),
      .datain(data0_i), .src_rdy_i(src0_rdy_i), .dst_rdy_o(dst0_rdy_o),
      .dataout(data0_int), .src_rdy_o(src0_rdy_int), .dst_rdy_i(dst0_rdy_int));

   fifo_short #(.WIDTH(36)) mux_fifo_in1
     (.clk(clk), .reset(reset), .clear(clear),
      .datain(data1_i), .src_rdy_i(src1_rdy_i), .dst_rdy_o(dst1_rdy_o),
      .dataout(data1_int), .src_rdy_o(src1_rdy_int), .dst_rdy_i(dst1_rdy_int));

   fifo_short #(.WIDTH(36)) mux_fifo_in2
     (.clk(clk), .reset(reset), .clear(clear),
      .datain(data2_i), .src_rdy_i(src2_rdy_i), .dst_rdy_o(dst2_rdy_o),
      .dataout(data2_int), .src_rdy_o(src2_rdy_int), .dst_rdy_i(dst2_rdy_int));

   localparam MUX_IDLE0 = 0;
   localparam MUX_DATA0 = 1;
   localparam MUX_IDLE1 = 2;
   localparam MUX_DATA1 = 3;
   localparam MUX_IDLE2 = 4;
   localparam MUX_DATA2 = 5;
   
   reg [2:0] 	  state;

   wire 	  eof0 = data0_int[33];
   wire 	  eof1 = data1_int[33];
   wire 	  eof2 = data2_int[33];
   
   wire [35:0] 	  data_int;
   wire 	  src_rdy_int, dst_rdy_int;
   
   // wtf?
   always @(posedge clk)
     if(reset | clear)
       state <= MUX_IDLE0;
     else
       case(state)
	 MUX_IDLE0 :
	   if(src0_rdy_int)
	     state <= MUX_DATA0;
	   else if(src1_rdy_int)
	     state <= MUX_DATA1;

	 MUX_DATA0 :
	   if(src0_rdy_int & dst_rdy_int & eof0)
	     state <= MUX_IDLE1;

	 MUX_IDLE1 :
	   if(src1_rdy_int)
	     state <= MUX_DATA1;
	   else if(src2_rdy_int)
	     state <= MUX_DATA2;
	   
	 MUX_DATA1 :
	   if(src1_rdy_int & dst_rdy_int & eof1)
	     state <= MUX_IDLE2;
       
	 MUX_IDLE2 :
	   if(src2_rdy_int)
	     state <= MUX_DATA2;
	   else if(src0_rdy_int)
	     state <= MUX_DATA0;
	   
	 MUX_DATA2 :
	   if(src1_rdy_int & dst_rdy_int & eof2)
	     state <= MUX_IDLE0;
	 
	 default :
	   state <= MUX_IDLE0;
       endcase // case (state)

   assign dst0_rdy_int = (state==MUX_DATA0) ? dst_rdy_int : 0;
   assign dst1_rdy_int = (state==MUX_DATA1) ? dst_rdy_int : 0;
   assign dst2_rdy_int = (state==MUX_DATA2) ? dst_rdy_int : 0;
   assign src_rdy_int = (state==MUX_DATA0) ? src0_rdy_int : (state==MUX_DATA1) ? src1_rdy_int : (state== MUX_DATA2) ? src2_rdy_int : 0;
   assign data_int = (state==MUX_DATA0) ? data0_int : (state==MUX_DATA1) ? data1_int : data2_int;
   
   fifo_short #(.WIDTH(36)) mux_fifo
     (.clk(clk), .reset(reset), .clear(clear),
      .datain(data_int), .src_rdy_i(src_rdy_int), .dst_rdy_o(dst_rdy_int),
      .dataout(data_o), .src_rdy_o(src_rdy_o), .dst_rdy_i(dst_rdy_i));
endmodule // fifo36_demux
